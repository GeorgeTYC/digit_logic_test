module debounce(clk,key,key_out);
